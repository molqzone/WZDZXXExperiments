module top (
        input      clock,
        input      reset
    );



endmodule
